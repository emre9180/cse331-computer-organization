module and_32bit(input [31:0] input1, input [31:0] input2, output [31:0] s);

and and1(s[0], input1[0], input2[0]);
and and2(s[1], input1[1], input2[1]);
and and3(s[2], input1[2], input2[2]);
and and4(s[3], input1[3], input2[3]);
and and5(s[4], input1[4], input2[4]);
and and6(s[5], input1[5], input2[5]);
and and7(s[6], input1[6], input2[6]);
and and8(s[7], input1[7], input2[7]);
and and9(s[8], input1[8], input2[8]);
and and10(s[9], input1[9], input2[9]);
and and11(s[10], input1[10], input2[10]);
and and12(s[11], input1[11], input2[11]);
and and13(s[12], input1[12], input2[12]);
and and14(s[13], input1[13], input2[13]);
and and15(s[14], input1[14], input2[14]);
and and16(s[15], input1[15], input2[15]);
and and17(s[16], input1[16], input2[16]);
and and18(s[17], input1[17], input2[17]);
and and19(s[18], input1[18], input2[18]);
and and20(s[19], input1[19], input2[19]);
and and21(s[20], input1[20], input2[20]);
and and22(s[21], input1[21], input2[21]);
and and223(s[22], input1[22], input2[22]);
and and24(s[23], input1[23], input2[23]);
and and25(s[24], input1[24], input2[24]);
and and26(s[25], input1[25], input2[25]);
and and27(s[26], input1[26], input2[26]);
and and28(s[27], input1[27], input2[27]);
and and29(s[28], input1[28], input2[28]);
and and30(s[29], input1[29], input2[29]);
and and31(s[30], input1[30], input2[30]);
and and32(s[31], input1[31], input2[31]);

endmodule
