module xor_32bit(input [31:0] input1, input [31:0] input2, output [31:0] s);

xor xor1(s[0], input1[0], input2[0]);
xor xor2(s[1], input1[1], input2[1]);
xor xor3(s[2], input1[2], input2[2]);
xor xor4(s[3], input1[3], input2[3]);
xor xor5(s[4], input1[4], input2[4]);
xor xor6(s[5], input1[5], input2[5]);
xor xor7(s[6], input1[6], input2[6]);
xor xor8(s[7], input1[7], input2[7]);
xor xor9(s[8], input1[8], input2[8]);
xor xor10(s[9], input1[9], input2[9]);
xor xor11(s[10], input1[10], input2[10]);
xor xor12(s[11], input1[11], input2[11]);
xor xor13(s[12], input1[12], input2[12]);
xor xor14(s[13], input1[13], input2[13]);
xor xor15(s[14], input1[14], input2[14]);
xor xor16(s[15], input1[15], input2[15]);
xor xor17(s[16], input1[16], input2[16]);
xor xor18(s[17], input1[17], input2[17]);
xor xor19(s[18], input1[18], input2[18]);
xor xor20(s[19], input1[19], input2[19]);
xor xor21(s[20], input1[20], input2[20]);
xor xor22(s[21], input1[21], input2[21]);
xor xor23(s[22], input1[22], input2[22]);
xor xor24(s[23], input1[23], input2[23]);
xor xor25(s[24], input1[24], input2[24]);
xor xor26(s[25], input1[25], input2[25]);
xor xor27(s[26], input1[26], input2[26]);
xor xor28(s[27], input1[27], input2[27]);
xor xor29(s[28], input1[28], input2[28]);
xor xor30(s[29], input1[29], input2[29]);
xor xor31(s[30], input1[30], input2[30]);
xor xor32(s[31], input1[31], input2[31]);

endmodule
