module and_16bit(input [15:0] input1, input [15:0] input2, output [15:0] s);

and and1(s[0], input1[0], input2[0]);
and and2(s[1], input1[1], input2[1]);
and and3(s[2], input1[2], input2[2]);
and and4(s[3], input1[3], input2[3]);
and and5(s[4], input1[4], input2[4]);
and and6(s[5], input1[5], input2[5]);
and and7(s[6], input1[6], input2[6]);
and and8(s[7], input1[7], input2[7]);
and and9(s[8], input1[8], input2[8]);
and and10(s[9], input1[9], input2[9]);
and and11(s[10], input1[10], input2[10]);
and and12(s[11], input1[11], input2[11]);
and and13(s[12], input1[12], input2[12]);
and and14(s[13], input1[13], input2[13]);
and and15(s[14], input1[14], input2[14]);
and and16(s[15], input1[15], input2[15]);


endmodule
