module or_32bit(input [31:0] input1, input [31:0] input2, output [31:0] s);

or or1(s[0], input1[0], input2[0]);
or or2(s[1], input1[1], input2[1]);
or or3(s[2], input1[2], input2[2]);
or or4(s[3], input1[3], input2[3]);
or or5(s[4], input1[4], input2[4]);
or or6(s[5], input1[5], input2[5]);
or or7(s[6], input1[6], input2[6]);
or or8(s[7], input1[7], input2[7]);
or or9(s[8], input1[8], input2[8]);
or or10(s[9], input1[9], input2[9]);
or or11(s[10], input1[10], input2[10]);
or or12(s[11], input1[11], input2[11]);
or or13(s[12], input1[12], input2[12]);
or or14(s[13], input1[13], input2[13]);
or or15(s[14], input1[14], input2[14]);
or or16(s[15], input1[15], input2[15]);
or or17(s[16], input1[16], input2[16]);
or or18(s[17], input1[17], input2[17]);
or or19(s[18], input1[18], input2[18]);
or or20(s[19], input1[19], input2[19]);
or or21(s[20], input1[20], input2[20]);
or or22(s[21], input1[21], input2[21]);
or or23(s[22], input1[22], input2[22]);
or or24(s[23], input1[23], input2[23]);
or or25(s[24], input1[24], input2[24]);
or or26(s[25], input1[25], input2[25]);
or or27(s[26], input1[26], input2[26]);
or or28(s[27], input1[27], input2[27]);
or or29(s[28], input1[28], input2[28]);
or or30(s[29], input1[29], input2[29]);
or or31(s[30], input1[30], input2[30]);
or or32(s[31], input1[31], input2[31]);

endmodule
