module not_32bit(input [31:0] input1, output [31:0] result);

not not1(result[0], input1[0]);
not not2(result[1], input1[1]);
not not3(result[2], input1[2]);
not not4(result[3], input1[3]);
not not5(result[4], input1[4]);
not not6(result[5], input1[5]);
not not7(result[6], input1[6]);
not not8(result[7], input1[7]);
not not9(result[8], input1[8]);
not not10(result[9], input1[9]);
not not11(result[10], input1[10]);
not not12(result[11], input1[11]);
not not13(result[12], input1[12]);
not not14(result[13], input1[13]);
not not15(result[14], input1[14]);
not not16(result[15], input1[15]);
not not17(result[16], input1[16]);
not not18(result[17], input1[17]);
not not19(result[18], input1[18]);
not not20(result[19], input1[19]);
not not21(result[20], input1[20]);
not not22(result[21], input1[21]);
not not23(result[22], input1[22]);
not not24(result[23], input1[23]);
not not25(result[24], input1[24]);
not not26(result[25], input1[25]);
not not27(result[26], input1[26]);
not not28(result[27], input1[27]);
not not29(result[28], input1[28]);
not not30(result[29], input1[29]);
not not31(result[30], input1[30]);
not not32(result[31], input1[31]);

endmodule